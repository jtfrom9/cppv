module test();
   initial begin
      $display("hello, test.v");
   end
endmodule

     
